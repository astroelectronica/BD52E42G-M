.title KiCad schematic
.include "C:/AE/BD52E42G/models/BD52E42G.lib"
.include "C:/AE/BD52E42G/models/C2012C0G2W101J060AA_p.mod"
.include "C:/AE/BD52E42G/models/C2012JB2E102M085AA_p.mod"
.include "C:/AE/BD52E42G/models/C2012X7R2A104M125AA_p.mod"
R1 VDD /OUT {RPU}
V1 VDD 0 {VSUPPLY}
XU2 VDD 0 C2012X7R2A104M125AA_p
XU4 /OUT 0 C2012JB2E102M085AA_p
XU1 /OUT VDD 0 unconnected-_U1-PadNC_ /CT BD52E42G
XU3 /CT 0 C2012C0G2W101J060AA_p
.end
